module orgate(output o, input a,b);
    assign o = a | b;
endmodule
