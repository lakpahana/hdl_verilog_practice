module andgate (output o, input a, input b);
  assign o = a & b;
endmodule
